'timescale 1ms/10ns
mdoule t05_SPI_tb; 