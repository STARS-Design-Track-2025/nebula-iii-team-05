// `timescale 1ms/10ps

typedef enum logic [2:0] {
    LEFT=0,
    RIGHT,
    TRACK,
    BACKTRACK,
    FINISH,
    INIT,
    SEND
} state_cb;

module t05_cb_synthesis_tb;
    logic clk, reset, char_found;
    logic [3:0] finished;
    logic [6:0] max_index;
    logic [70:0] h_element;
    //logic [2:0] curr_process;
    logic [127:0] char_path;
    logic [7:0] char_index;
    logic [6:0] curr_index;
    state_cb state;
    logic [70:0] htree [127:0];
    logic [127:0] curr_path;
    logic [8:0] least1;
    logic [8:0] least2;
    logic [8:0] header;
    logic [6:0] track_length;
    logic [6:0] pos;
    logic mid_reset;
    logic [7:0] count;
    logic enable;
    logic bit1;
    logic write_finish;
    logic wait_cycle;

    always #5 clk = ~clk;
    t05_cb_synthesis cb1(.clk(clk), .write_finish(write_finish), .track_length(track_length), .pos(pos), .least1(least1), .least2(least2), .rst(reset), .max_index(max_index), .curr_path(curr_path), .curr_index(curr_index), .h_element(h_element), .curr_state(state), .char_path(char_path), .char_index(char_index), .char_found(char_found), .finished(finished), .wait_cycle(wait_cycle));
    t05_header_synthesis hd1 (.clk(clk), .write_finish(write_finish), .rst(reset), .bit1(bit1), .enable(enable), .char_index(char_index), .char_path(char_path), .char_found(char_found), .least1(least1), .least2(least2), .header(header));
    task reset_fsm();
      begin
        reset = 1;
        @(posedge clk);
        reset = 0;
        @(posedge clk);
      end
    endtask

//     task set_inputs(logic [6:0] max_index1, logic [70:0] h_element1);
//       begin
//         max_index = max_index1;
//         h_element = h_element1;
//         @(posedge clk);
//       end
//     endtask

//     initial begin
//       $dumpfile("t05_cb_synthesis.vcd"); //change the vcd vile name to your source file name
//       $dumpvars(0, t05_cb_synthesis_tb);
      
//       clk = 0;
//       reset = 0;
//       h_element = {{7'd8}, {1'b1, 8'd6}, {1'b1, 8'd7}, {46'd52}};
//       max_index = 8;
//       //header = 0;
//       htree[0] = {{7'd8}, {1'b0, 8'd67}, {1'b0, 8'd66}, {46'd5}}; // max_index=8, C=2, B=3, sum=5
//       htree[1] = {{7'd8}, {1'b0, 8'd68}, {1'b0, 8'd69}, {46'd7}}; // max_index=8, D=3, E=4, sum=7
//       htree[2] = {{7'd8}, {1'b0, 8'd72}, {1'b0, 8'd73}, {46'd8}}; // max_index=8, H=4, I=4, sum=8
//       htree[3] = {{7'd8}, {1'b1, 8'd0}, {1'b0, 8'd65}, {46'd10}}; // max_index=8, A=5, index0=5, sum=10
//       htree[4] = {{7'd8}, {1'b0, 8'd70}, {1'b1, 8'd1}, {46'd13}}; // max_index=8, F=6, index1=7, sum=13
//       htree[5] = {{7'd8}, {1'b0, 8'd71}, {1'b1, 8'd2}, {46'd15}}; // max_index=8, G=7, index2=8, sum=15
//       htree[6] = {{7'd8}, {1'b1, 8'd3}, {1'b1, 8'd4}, {46'd23}}; // max_index=8, index3=10, index4=13, sum=23
//       htree[7] = {{7'd8}, {1'b0, 8'd74}, {1'b1, 8'd5}, {46'd29}}; // max_index=8, J=14, index5=15, sum=29
//       htree[8] = {{7'd8}, {1'b1, 8'd6}, {1'b1, 8'd7}, {46'd52}}; // max_index=8, index6=23, index7=29, sum=52
      
//       reset_fsm();
//       $display("STATE: %d", state);
//       set_inputs(8, htree[8]); 
//       $display("STATE: %d", state);
//       //@(posedge clk);
//       set_inputs(8, htree[curr_index]);
//       $display("STATE: %d", state);
//       //@(posedge clk);
//       set_inputs(8, htree[curr_index]);
//       $display("STATE: %d", state); 
//       //@(posedge clk);
//       set_inputs(8, htree[curr_index]);
//       $display("STATE: %d", state); 
//       //@(posedge clk);
//       set_inputs(8, htree[curr_index]);
//       $display("STATE: %d", state); 
//       //@(posedge clk);
//       set_inputs(8, htree[curr_index]);
//       $display("STATE: %d", state); 
//       //@(posedge clk);
//       set_inputs(8, htree[curr_index]);
//       $display("STATE: %d", state); 
//       //@(posedge clk);
//       set_inputs(8, htree[curr_index]);
//       $display("STATE: %d", state); 
//       //@(posedge clk);
//       set_inputs(8, htree[curr_index]);
//       $display("STATE: %d", state);  
//       //@(posedge clk);
//       set_inputs(8, htree[curr_index]);
//       $display("STATE: %d", state);
//       //@(posedge clk);
//       set_inputs(8, htree[curr_index]);
//       $display("STATE: %d", state);
//       //@(posedge clk);
//       set_inputs(8, htree[curr_index]);
//       $display("STATE: %d", state); 
//       //@(posedge clk);
//       set_inputs(8, htree[curr_index]);
//       $display("STATE: %d", state); 
//       //@(posedge clk);
//       set_inputs(8, htree[curr_index]);
//       $display("STATE: %d", state); 
//       //@(posedge clk);
//       set_inputs(8, htree[curr_index]);
//       $display("STATE: %d", state); 
//       //@(posedge clk);
//       set_inputs(8, htree[curr_index]);
//       $display("STATE: %d", state); 
//       //@(posedge clk);
//       set_inputs(8, htree[curr_index]);
//       $display("STATE: %d", state); 
//       //@(posedge clk);
//       set_inputs(8, htree[curr_index]);
//       $display("STATE: %d", state);  
//       //@(posedge clk);
//       set_inputs(8, htree[curr_index]);
//       $display("STATE: %d", state); 
//       //@(posedge clk);
//       set_inputs(8, htree[curr_index]);
//       $display("STATE: %d", state); 
//       //@(posedge clk);
//       set_inputs(8, htree[curr_index]);
//       $display("STATE: %d", state); 
//       //@(posedge clk);
//       set_inputs(8, htree[curr_index]);
//       $display("STATE: %d", state); 
//       //@(posedge clk);
//       set_inputs(8, htree[curr_index]);
//       $display("STATE: %d", state); 
//       //@(posedge clk);
//       set_inputs(8, htree[curr_index]);
//       $display("STATE: %d", state); 
//       //@(posedge clk);
//       set_inputs(8, htree[curr_index]);
//       $display("STATE: %d", state); 
//       //@(posedge clk);
//       set_inputs(8, htree[curr_index]);
//       $display("STATE: %d", state);  
//       //@(posedge clk);
//       set_inputs(8, htree[curr_index]);
//       $display("STATE: %d", state); 
//       //@(posedge clk);
//       set_inputs(8, htree[curr_index]);
//       $display("STATE: %d", state); 
//       //@(posedge clk);
//       set_inputs(8, htree[curr_index]);
//       $display("STATE: %d", state); 
//       //@(posedge clk);
//       set_inputs(8, htree[curr_index]);
//       $display("STATE: %d", state); 
//       //@(posedge clk);
//       set_inputs(8, htree[curr_index]);
//       $display("STATE: %d", state); 
//       //@(posedge clk);
//       set_inputs(8, htree[curr_index]);
//       $display("STATE: %d", state); 
//       //@(posedge clk);
//       set_inputs(8, htree[curr_index]);
//       $display("STATE: %d", state); 
//       //@(posedge clk);
//       set_inputs(8, htree[curr_index]);
//       $display("STATE: %d", state);  
//       //@(posedge clk);
//       set_inputs(8, htree[curr_index]);
//       $display("STATE: %d", state); 
//       $display("STATE: %d", state);
//       //@(posedge clk);
//       set_inputs(8, htree[curr_index]);
//       $display("STATE: %d", state);
//       //@(posedge clk);
//       set_inputs(8, htree[curr_index]);
//       $display("STATE: %d", state); 
//       //@(posedge clk);
//       set_inputs(8, htree[curr_index]);
//       $display("STATE: %d", state); 
//       //@(posedge clk);
//       set_inputs(8, htree[curr_index]);
//       $display("STATE: %d", state); 
//       //@(posedge clk);
//       set_inputs(8, htree[curr_index]);
//       $display("STATE: %d", state); 
//       //@(posedge clk);
//       set_inputs(8, htree[curr_index]);
//       $display("STATE: %d", state); 
//       //@(posedge clk);
//       set_inputs(8, htree[curr_index]);
//       $display("STATE: %d", state); 
//       //@(posedge clk);
//       set_inputs(8, htree[curr_index]);
//       $display("STATE: %d", state);  
//       //@(posedge clk);
//       set_inputs(8, htree[curr_index]);
//       $display("STATE: %d", state);
//       //@(posedge clk);
//       set_inputs(8, htree[curr_index]);
//       $display("STATE: %d", state);
//       //@(posedge clk);
//       set_inputs(8, htree[curr_index]);
//       $display("STATE: %d", state); 
//       //@(posedge clk);
//       set_inputs(8, htree[curr_index]);
//       $display("STATE: %d", state); 
//       //@(posedge clk);
//       set_inputs(8, htree[curr_index]);
//       $display("STATE: %d", state); 
//       //@(posedge clk);
//       set_inputs(8, htree[curr_index]);
//       $display("STATE: %d", state); 
//       //@(posedge clk);
//       set_inputs(8, htree[curr_index]);
//       $display("STATE: %d", state); 
//       //@(posedge clk);
//       set_inputs(8, htree[curr_index]);
//       $display("STATE: %d", state); 
//       //@(posedge clk);
//       set_inputs(8, htree[curr_index]);
//       $display("STATE: %d", state);  
//       //@(posedge clk);
//       set_inputs(8, htree[curr_index]);
//       $display("STATE: %d", state); 
//       //@(posedge clk);
//       set_inputs(8, htree[curr_index]);
//       $display("STATE: %d", state); 
//       //@(posedge clk);
//       set_inputs(8, htree[curr_index]);
//       $display("STATE: %d", state); 
//       //@(posedge clk);
//       set_inputs(8, htree[curr_index]);
//       $display("STATE: %d", state); 
//       //@(posedge clk);
//       set_inputs(8, htree[curr_index]);
//       $display("STATE: %d", state); 
//       //@(posedge clk);
//       set_inputs(8, htree[curr_index]);
//       $display("STATE: %d", state); 
//       set_inputs(8, htree[curr_index]);
//       $display("STATE: %d", state);
//       //@(posedge clk);
//       set_inputs(8, htree[curr_index]);
//       $display("STATE: %d", state); 
//       //@(posedge clk);
//       set_inputs(8, htree[curr_index]);
//       $display("STATE: %d", state); 
//       //@(posedge clk);
//       set_inputs(8, htree[curr_index]);
//       $display("STATE: %d", state); 
//       //@(posedge clk);
//       set_inputs(8, htree[curr_index]);
//       $display("STATE: %d", state); 
//       //@(posedge clk);
//       set_inputs(8, htree[curr_index]);
//       $display("STATE: %d", state); 
//       //@(posedge clk);
//       set_inputs(8, htree[curr_index]);
//       $display("STATE: %d", state); 
//       //@(posedge clk);
//       set_inputs(8, htree[curr_index]);
//       $display("STATE: %d", state);  
//       //@(posedge clk);
//       set_inputs(8, htree[curr_index]);
//       $display("STATE: %d", state); 
//       //@(posedge clk);
//       set_inputs(8, htree[curr_index]);
//       $display("STATE: %d", state); 
//       //@(posedge clk);
//       set_inputs(8, htree[curr_index]);
//       $display("STATE: %d", state); 
//       //@(posedge clk);
//       set_inputs(8, htree[curr_index]);
//       $display("STATE: %d", state); 
//       //@(posedge clk);
//       set_inputs(8, htree[curr_index]);
//       $display("STATE: %d", state); 
//       //@(posedge clk);
//       set_inputs(8, htree[curr_index]);
//       $display("STATE: %d", state); 
//       set_inputs(8, htree[curr_index]);
//       $display("STATE: %d", state);
//       //@(posedge clk);
//       set_inputs(8, htree[curr_index]);
//       $display("STATE: %d", state); 
//       //@(posedge clk);
//       set_inputs(8, htree[curr_index]);
//       $display("STATE: %d", state); 
//       //@(posedge clk);
//       set_inputs(8, htree[curr_index]);
//       $display("STATE: %d", state); 
//       //@(posedge clk);
//       set_inputs(8, htree[curr_index]);
//       $display("STATE: %d", state); 
//       //@(posedge clk);
//       set_inputs(8, htree[curr_index]);
//       $display("STATE: %d", state); 
//       //@(posedge clk);
//       set_inputs(8, htree[curr_index]);
//       $display("STATE: %d", state); 
//       //@(posedge clk);
//       set_inputs(8, htree[curr_index]);
//       $display("STATE: %d", state);  
//       //@(posedge clk);
//       set_inputs(8, htree[curr_index]);
//       $display("STATE: %d", state); 
//       //@(posedge clk);
//       set_inputs(8, htree[curr_index]);
//       $display("STATE: %d", state); 
//       //@(posedge clk);
//       set_inputs(8, htree[curr_index]);
//       $display("STATE: %d", state); 
//       //@(posedge clk);
//       set_inputs(8, htree[curr_index]);
//       $display("STATE: %d", state); 
//       //@(posedge clk);
//       set_inputs(8, htree[curr_index]);
//       $display("STATE: %d", state); 
//       //@(posedge clk);
//       set_inputs(8, htree[curr_index]);
//       $display("STATE: %d", state); 
//       set_inputs(8, htree[curr_index]);
//       $display("STATE: %d", state);
//       //@(posedge clk);
//       set_inputs(8, htree[curr_index]);
//       $display("STATE: %d", state); 
//       //@(posedge clk);
//       set_inputs(8, htree[curr_index]);
//       $display("STATE: %d", state); 
//       //@(posedge clk);
//       set_inputs(8, htree[curr_index]);
//       $display("STATE: %d", state); 
//       //@(posedge clk);
//       set_inputs(8, htree[curr_index]);
//       $display("STATE: %d", state); 
//       //@(posedge clk);
//       set_inputs(8, htree[curr_index]);
//       $display("STATE: %d", state); 
//       //@(posedge clk);
//       set_inputs(8, htree[curr_index]);
//       $display("STATE: %d", state); 
//       //@(posedge clk);
//       set_inputs(8, htree[curr_index]);
//       $display("STATE: %d", state);  
//       //@(posedge clk);
//       set_inputs(8, htree[curr_index]);
//       $display("STATE: %d", state); 
//       //@(posedge clk);
//       set_inputs(8, htree[curr_index]);
//       $display("STATE: %d", state); 
//       //@(posedge clk);
//       set_inputs(8, htree[curr_index]);
//       $display("STATE: %d", state); 
//       //@(posedge clk);
//       set_inputs(8, htree[curr_index]);
//       $display("STATE: %d", state); 
//       //@(posedge clk);
//       set_inputs(8, htree[curr_index]);
//       $display("STATE: %d", state); 
//       //@(posedge clk);
//       set_inputs(8, htree[curr_index]);
//       $display("STATE: %d", state); 
//       set_inputs(8, htree[curr_index]);
//       $display("STATE: %d", state);
//       //@(posedge clk);
//       set_inputs(8, htree[curr_index]);
//       $display("STATE: %d", state); 
//       //@(posedge clk);
//       set_inputs(8, htree[curr_index]);
//       $display("STATE: %d", state); 
//       //@(posedge clk);
//       set_inputs(8, htree[curr_index]);
//       $display("STATE: %d", state); 
//       //@(posedge clk);
//       set_inputs(8, htree[curr_index]);
//       $display("STATE: %d", state); 
//       //@(posedge clk);
//       set_inputs(8, htree[curr_index]);
//       $display("STATE: %d", state); 
//       //@(posedge clk);
//       set_inputs(8, htree[curr_index]);
//       $display("STATE: %d", state); 
//       //@(posedge clk);
//       set_inputs(8, htree[curr_index]);
//       $display("STATE: %d", state);  
//       //@(posedge clk);
//       set_inputs(8, htree[curr_index]);
//       $display("STATE: %d", state); 
//       //@(posedge clk);
//       set_inputs(8, htree[curr_index]);
//       $display("STATE: %d", state); 
//       //@(posedge clk);
//       set_inputs(8, htree[curr_index]);
//       $display("STATE: %d", state); 
//       //@(posedge clk);
//       set_inputs(8, htree[curr_index]);
//       $display("STATE: %d", state); 
//       //@(posedge clk);
//       set_inputs(8, htree[curr_index]);
//       $display("STATE: %d", state); 
//       //@(posedge clk);
//       set_inputs(8, htree[curr_index]);
//       $display("STATE: %d", state); 

      #10;

//       #1 $finish;

//     end
  
// endmodule
  