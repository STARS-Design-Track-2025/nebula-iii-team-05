`timescale 1ms/10ps

typedef enum logic [3:0] {
    INIT, // initial (set if enable for the hd_decode module isn't high)
    READ_NUM_LEFTS, // reads the 9 bit chunk of the number of lefts after moving right for the left char stored in the header
    READ_LEADING_BIT, // read leading bit checks if there is a backtrack (0) or if another char was found (1)
    READ_CHAR, // read 8 bits of the char from data_in after reading the leading bit(s)
    UPDATE_PATH, // after getting the character, use the # of backtrack and the bit after the char to update the path
    WRITE_PATH, // once a full path is found, (after a char was found and corresponding path was updated with correct digits), send the path to SRAM with the curr char index
    READ_TOT_CHAR, // read the total number chars in the file after the whole binary tree was turned into a codebook  
    FINISH // finished writing all char codes from header
} state_hd;

module t05_hd_decode_tb;
    logic clk, reset;
    logic hd_enable;
    logic [7:0] SPI_data_in; // read byte of header from SPI
    logic read_en_SPI;
    logic [127:0] SRAM_data_out; // write a char path to SRAM
    logic SRAM_write_en;
    logic [935:0] SPI_data_arr; // enough for 256 characters and an average of 2 zeroes per char
    logic [31:0] tot_chars;
    logic finished;

    always #5 clk = ~clk;
    t05_hd_decode hd1 (.clk(clk), .rst(reset), .finished(finished), .tot_chars(tot_chars), .hd_enable(1'b1), .SPI_data_in(SPI_data_in), .SPI_read_en(read_en_SPI), .SRAM_data_out(SRAM_data_out), .SRAM_write_en(SRAM_write_en));
    task reset_fsm();
      begin
        reset = 1;
        @(posedge clk);
        reset = 0;
        @(posedge clk);
      end
    endtask

    task set_inputs(logic [7:0] SPI_data, logic SPI_enable);
      begin
        //if (SPI_enable) begin
            SPI_data_in = SPI_data;
            @(posedge clk);
        //end
      end
    endtask

    task automatic feed_spi_stream(input logic [935:0] spi_data, input int num_bytes);
    //SPI_data_in = spi_data[263-: 8];
    //int i = 0;
      //while (!finished) begin
      for (int i = 0; i < 117; i++) begin
        @(posedge clk);
        while (!read_en_SPI) @(posedge clk);

        SPI_data_in = spi_data[935 - 8*i -: 8];
        //i++;
        @(posedge clk);
    end
endtask

    initial begin
      $dumpfile("t05_hd_decode.vcd"); //change the vcd vile name to your source file name
      $dumpvars(0, t05_hd_decode_tb);
      
      clk = 0;
      reset = 0;
      //SPI_data_arr[263:0] = 264'b0;
      //SPI_data_arr[263:0] = {{1'b1, 8'd67, 9'b100000100}, {1'b1, 8'd66, 1'b0}, + {1'b1, 8'd65, 1'b0}, {1'b1, 8'd70, 9'b100000001}, {1'b1, 8'd71, 2'b0}, {1'b1, 8'd74, 9'b100000001}, {1'b1, 8'd68, 9'b100000011},{1'b1, 8'd69, 1'b0}, {1'b1, 8'd75, 1'b0}, {1'b1, 8'd72, 9'b100000001}, {1'b1, 8'd73, 4'b0}, {1'b1, 8'b00001010}, {32'd11}, {69'b0}};
      
      //LONG HTREE
      // SPI_data_arr[911:0] = {880'b101011110100000001101011101100000001101011100100000001101011011100000001101011010100000001101011001100000001101011000100000001101010111100000001101010110100000001101010101100000001101010100100000001101010011100000001101010010100000001101010001100000001101010000100000001101011110100000001101011101100000001101011100100000001101011011100000001101011010100000001101011001100000001101011000100000001101010111100000001101010110100000001101010101100000001101010100100000001101010011100000001101010010100000001101010001100000001101010000100000001101001111100000001101001110100000001101001101100000001101001100100000001101001011100000001101001010100000001101001001100000001101001000100000001101000111100000001101000110100000001101000101100000001101000100100000001101000011100000001101000010100000001101000001100000001100000000100000001100000001000000000000000000000000000100001010, 32'd666};
      // reset_fsm();
      // feed_spi_stream(SPI_data_arr, 114);
      
      SPI_data_arr[935:0] = {904'b1011011111000001011001011100101110000100000001100101111001011100011000000101001100000101110010100000001100110001000101110011100000011100110010010111010010000000110011001100101110101100000010100110100010110111110000010110010111001011100001000000011001011110010111000110000001010011000001011100101000000011001100010001011100111000000111001100100101110100100000001100110011001011101011000000101001101000101110110100000001100110101000010101111110000010110001111001011000001000000011000111110010110000110000001010010000001011000101000000011001000010001011000111000000111001000100101100100100000001100100011001011001011000000101001001000101100110100000001100100101000010110011110000010010010011001011010001000000011001001110010110100110000001010010100001011010101000000011001010010001011010111000000111001010100101101100100000001100101011001011011011000000101001011000101101110100000001100101101000000100001010, 32'd2626};
      reset_fsm();
      feed_spi_stream(SPI_data_arr, 117);
      // SPI_data_arr[263:0] = {128'b10000, {1'b1, 8'd67}, {1'b1, 8'd66, 1'b0}, + {1'b1, 8'd65, 1'b0}, {1'b1, 8'd70}, {1'b1, 8'd71, 2'b0}, {1'b1, 8'd74}, {1'b1, 8'd68}, {1'b1, 8'd75}, {1'b1, 8'd69, 1'b0}, {1'b1, 8'd72}, {1'b1, 8'd73, 4'b0}, {32'd10}, {12'b0}};
//       set_inputs(SPI_data_arr[263:256], read_en_SPI);
//       while (!read_en_SPI) begin
//         set_inputs(SPI_data_arr[263:256], read_en_SPI);
//       end
//       set_inputs(SPI_data_arr[255:248], read_en_SPI);
//       while (!read_en_SPI) begin
//         set_inputs(SPI_data_arr[255:248], read_en_SPI);
//       end
//        set_inputs(SPI_data_arr[247:240], read_en_SPI);
//       while (!read_en_SPI) begin
//         set_inputs(SPI_data_arr[247:240], read_en_SPI);
//       end
//       set_inputs(SPI_data_arr[239:232], read_en_SPI);
//       while (!read_en_SPI) begin
//         set_inputs(SPI_data_arr[239:232], read_en_SPI);
//       end
//       set_inputs(SPI_data_arr[231:224], read_en_SPI);
//       while (!read_en_SPI) begin
//         set_inputs(SPI_data_arr[231:224], read_en_SPI);
//       end
//       set_inputs(SPI_data_arr[223:216], read_en_SPI);
//       while (!read_en_SPI) begin
//         set_inputs(SPI_data_arr[223:216], read_en_SPI);
//       end
//       set_inputs(SPI_data_arr[215:208], read_en_SPI);
//       while (!read_en_SPI) begin
//       set_inputs(SPI_data_arr[215:208], read_en_SPI);
//       end

//       set_inputs(SPI_data_arr[207:200], read_en_SPI);
//     while (!read_en_SPI) begin
//       set_inputs(SPI_data_arr[207:200], read_en_SPI);
//     end

    
//       set_inputs(SPI_data_arr[199:192], read_en_SPI);
//     while (!read_en_SPI) begin
//       set_inputs(SPI_data_arr[199:192], read_en_SPI);
//     end

//       set_inputs(SPI_data_arr[191:184], read_en_SPI);
//     while (!read_en_SPI) begin
//       set_inputs(SPI_data_arr[191:184], read_en_SPI);
//     end

//       set_inputs(SPI_data_arr[183:176], read_en_SPI);
//     while (!read_en_SPI) begin
//       set_inputs(SPI_data_arr[183:176], read_en_SPI);
//     end

//       set_inputs(SPI_data_arr[175:168], read_en_SPI);
//     while (!read_en_SPI) begin
//       set_inputs(SPI_data_arr[175:168], read_en_SPI);
//     end

//       set_inputs(SPI_data_arr[167:160], read_en_SPI);
//     while (!read_en_SPI) begin
//       set_inputs(SPI_data_arr[167:160], read_en_SPI);
//     end

//       set_inputs(SPI_data_arr[159:152], read_en_SPI);
//     while (!read_en_SPI) begin
//       set_inputs(SPI_data_arr[159:152], read_en_SPI);
//     end

//       set_inputs(SPI_data_arr[151:144], read_en_SPI);
//     while (!read_en_SPI) begin
//       set_inputs(SPI_data_arr[151:144], read_en_SPI);
//     end

//       set_inputs(SPI_data_arr[143:136], read_en_SPI);
//     while (!read_en_SPI) begin
//       set_inputs(SPI_data_arr[143:136], read_en_SPI);
//     end

//       set_inputs(SPI_data_arr[135:128], read_en_SPI);
//     while (!read_en_SPI) begin
//       set_inputs(SPI_data_arr[135:128], read_en_SPI);
//     end

//       set_inputs(SPI_data_arr[127:120], read_en_SPI);
//     while (!read_en_SPI) begin
//       set_inputs(SPI_data_arr[127:120], read_en_SPI);
//     end

//       set_inputs(SPI_data_arr[119:112], read_en_SPI);
//     while (!read_en_SPI) begin
//       set_inputs(SPI_data_arr[119:112], read_en_SPI);
//     end

//       set_inputs(SPI_data_arr[111:104], read_en_SPI);
//     while (!read_en_SPI) begin
//       set_inputs(SPI_data_arr[111:104], read_en_SPI);
//     end
      
//       set_inputs(SPI_data_arr[103:96], read_en_SPI);
//     while (!read_en_SPI) begin
//       set_inputs(SPI_data_arr[103:96], read_en_SPI);
//     end

//       set_inputs(SPI_data_arr[95:88], read_en_SPI);
//     while (!read_en_SPI) begin
//       set_inputs(SPI_data_arr[95:88], read_en_SPI);
//     end

//       set_inputs(SPI_data_arr[87:80], read_en_SPI);
//     while (!read_en_SPI) begin
//       set_inputs(SPI_data_arr[87:80], read_en_SPI);
//     end

//       set_inputs(SPI_data_arr[79:72], read_en_SPI);
//     while (!read_en_SPI) begin
//       set_inputs(SPI_data_arr[79:72], read_en_SPI);
//     end

//       set_inputs(SPI_data_arr[71:64], read_en_SPI);
//     while (!read_en_SPI) begin
//       set_inputs(SPI_data_arr[71:64], read_en_SPI);
//     end

//       set_inputs(SPI_data_arr[63:56], read_en_SPI);
//     while (!read_en_SPI) begin
//       set_inputs(SPI_data_arr[63:56], read_en_SPI);
//     end

//       set_inputs(SPI_data_arr[55:48], read_en_SPI);
//     while (!read_en_SPI) begin
//       set_inputs(SPI_data_arr[55:48], read_en_SPI);
//     end

//       set_inputs(SPI_data_arr[47:40], read_en_SPI);
//     while (!read_en_SPI) begin
//       set_inputs(SPI_data_arr[47:40], read_en_SPI);
//     end
      
//       set_inputs(SPI_data_arr[39:32], read_en_SPI);
//      // #500
//     while (!read_en_SPI) begin
//       set_inputs(SPI_data_arr[39:32], read_en_SPI);
//     end

//       set_inputs(SPI_data_arr[31:24], read_en_SPI);
//     while (!read_en_SPI) begin
//       set_inputs(SPI_data_arr[31:24], read_en_SPI);
//     end
 
//       set_inputs(SPI_data_arr[23:16], read_en_SPI);
//     while (!read_en_SPI) begin
//       set_inputs(SPI_data_arr[23:16], read_en_SPI);
//     end

//       set_inputs(SPI_data_arr[15:8], read_en_SPI);
//     while (!read_en_SPI) begin
//       set_inputs(SPI_data_arr[15:8], read_en_SPI);
//     end

//       set_inputs(SPI_data_arr[7:0], read_en_SPI);
    // while (!read_en_SPI) begin
    //   set_inputs(SPI_data_arr[7:0], read_en_SPI);
    // end
    
      #100;

      #1 $finish;

    end
  
endmodule
